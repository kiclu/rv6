`ifdef __ICARUS__
    `define program_hex_path "test/c/default/default.hex"
    `define mem_final_path   "test/out/tb_hart_mem.hex"
    `define finish $finish
`else
    `define program_hex_path "../test/c/default/default.hex"
    `define mem_final_path   "../test/out/tb_hart_mem.hex"
    `define finish $stop
`endif

`include "../hdl/config.v"

`timescale 1ns/1ps
module tb_hart_fib();

    wire           [63:0] b_addr_i;
    reg  [`imem_line-1:0] b_data_i;
    wire                  b_rd_i;
    reg                   b_dv_i;

    wire           [63:0] b_addr;

    reg  [`dmem_line-1:0] b_data_in;
    wire                  b_rd;
    reg                   b_dv;

    wire [`dmem_line-1:0] b_data_out;
    wire                  b_wr;

    reg                   rst_n;
    reg                   clk;

    reg [7:0] rom [0:4095];
    reg [7:0] ram [0:32767];

    initial begin
        b_data_i  = `imem_line'bZ;
        b_dv_i    = 1'b0;

        b_data_in = `dmem_line'bZ;
        b_dv      = 1'b0;

        rst_n     = 1'b0;

        clk       = 1'b1;

        forever #10 clk = ~clk;
    end

    initial $readmemh(`program_hex_path, rom, 0);

    initial begin
        for(integer i = 0; i < 4096; ++i) begin
            if(rom[i] === 8'bxxxxxxxx) rom[i] = 8'b0;
        end
        for(integer i = 0; i < 32768; ++i) ram[i] = 8'b0;
    end

    initial begin
        #40
        rst_n = 1'b1;
        #10000
        $writememh(`mem_final_path, ram, 0);
        `finish();
    end

    always @(posedge clk) begin
        if(b_rd_i) begin
            #80
            for(integer i = 0; i < `imem_line/8; ++i) begin
                b_data_i[8*i +: 8] = rom[b_addr_i + i - 64'h80000000];
            end
            b_dv_i = 1;
            #20
            b_data_i = `imem_line'bZ;
            b_dv_i   = 0;
        end
        if(b_rd) begin
            #80
            for(integer i = 0; i < `dmem_line/8; ++i) begin
                b_data_in[8*i +: 8] = ram[b_addr + i];
            end
            b_dv = 1;
            #20
            b_data_in = `dmem_line'bZ;
            b_dv      = 0;
        end
        if(b_wr) begin
            for(integer i = 0; i < `dmem_line/8; ++i) begin
                ram[b_addr + i] = b_data_out[8*i +: 8];
            end
        end
    end

    hart dut(
        .b_addr_i(b_addr_i),
        .b_data_i(b_data_i),
        .b_rd_i(b_rd_i),
        .b_dv_i(b_dv_i),

        .b_addr(b_addr),

        .b_data_in(b_data_in),
        .b_rd(b_rd),
        .b_dv(b_dv),

        .b_data_out(b_data_out),
        .b_wr(b_wr),

        .rst_n(rst_n),

        .clk(clk)
    );

endmodule
