/*
 * Copyright (C) 2023  Nikola Lukic <lukicn@protonmail.com>
 * This source describes Open Hardware and is licensed under the CERN-OHL-W v2
 *
 * You may redistribute and modify this documentation and make products
 * using it under the terms of the CERN-OHL-W v2 (https:/cern.ch/cern-ohl).
 * This documentation is distributed WITHOUT ANY EXPRESS OR IMPLIED
 * WARRANTY, INCLUDING OF MERCHANTABILITY, SATISFACTORY QUALITY
 * AND FITNESS FOR A PARTICULAR PURPOSE. Please see the CERN-OHL-W v2
 * for applicable conditions.
 *
 * Source location: https://www.github.com/kiclu/rv6
 *
 * As per CERN-OHL-W v2 section 4.1, should You produce hardware based on
 * these sources, You must maintain the Source Location visible on the
 * external case of any product you make using this documentation.
 */

module pd(
    input      [63:0] pc_in,
    input      [31:0] ir_in,

    output reg [63:0] pc_out,
    output reg [31:0] ir_out,

    input             stall,

    input             clk
);

    always @(negedge clk) begin
        if(!stall) begin
            casez(ir_in)
                default: begin
                    pc_out <= pc_in;
                    ir_out <= ir_in;
                end
            endcase
        end
    end

endmodule
